module top_module();
    
    reg [1:0] in;
    
    initial begin
    assign in = 2'b00;
    #10
    assign in = 2'b01;
    #10
    assign in = 2'b10;
    #10
    assign in = 2'b11;
    end
        
    wire out;
    andgate I0(.out(out), .in(in));
    
endmodule